typedef 8   NumInputs;
typedef 100 CyclesResolution;

typedef 8  NumLeds;
typedef 15 Log2LedPersistence;
typedef 7  Log2ErrorBlink;
